library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pck_definitions is
  constant num_bits : integer := 16;
  constant num_bits_int_part : integer := 4;
  constant num_bits_frac_part : integer := num_bits - num_bits_int_part;
  constant zero : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 0, num_bits );
  constant one : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4096, num_bits );
  constant a_to_1_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 64, num_bits );
  constant b_to_1_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 18143, num_bits );
  constant c_to_1_neg_expon : integer := 6;
  constant a_to_2_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 145, num_bits );
  constant b_to_2_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 14900, num_bits );
  constant c_to_2_neg_expon : integer := 5;
  constant a_to_3_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 20, num_bits );
  constant b_to_3_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 15942, num_bits );
  constant c_to_3_neg_expon : integer := 5;
  constant a_to_4_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -228, num_bits );
  constant b_to_4_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 17293, num_bits );
  constant c_to_4_neg_expon : integer := 5;
  constant a_to_5_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4324, num_bits );
  constant b_to_5_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -17293, num_bits );
  constant c_to_5_neg_expon : integer := 5;
  constant a_to_6_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4076, num_bits );
  constant b_to_6_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -15942, num_bits );
  constant c_to_6_neg_expon : integer := 5;
  constant a_to_7_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 3951, num_bits );
  constant b_to_7_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -14900, num_bits );
  constant c_to_7_neg_expon : integer := 5;
  constant a_to_8_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4032, num_bits );
  constant b_to_8_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -18143, num_bits );
  constant c_to_8_neg_expon : integer := 6;
  constant lambda_0 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -16384, num_bits );
  constant lambda_0_1_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -12288, num_bits );
  constant lambda_0_2_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -8192, num_bits );
  constant lambda_0_3_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -4096, num_bits );
  constant lambda_0_4_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 0, num_bits );
  constant lambda_0_5_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4096, num_bits );
  constant lambda_0_6_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 8192, num_bits );
  constant lambda_0_7_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 12288, num_bits );
  constant lambda_0_8_delta : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 16384, num_bits );
end package pck_definitions;
