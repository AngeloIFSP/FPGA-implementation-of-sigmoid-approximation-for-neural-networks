library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pck_definitions is
  constant num_bits : integer := 16;
  constant num_bits_int_part : integer := 4;
  constant num_bits_frac_part : integer := num_bits - num_bits_int_part;
  constant zero : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 0, num_bits );
  constant one : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4096, num_bits );
  constant limit_minus_8 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -32768, num_bits );
  constant limit_minus_4_5 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -18432, num_bits );
  constant limit_minus_3 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -12288, num_bits );
  constant limit_minus_2 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -8192, num_bits );
  constant limit_minus_1 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( -4096, num_bits );
  constant limit_plus_1 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4096, num_bits );
  constant limit_plus_2 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 8192, num_bits );
  constant limit_plus_3 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 12288, num_bits );
  constant limit_plus_4_5 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 18432, num_bits );
  constant limit_plus_8 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 32767, num_bits );
  constant coef_1 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 10, num_bits );
  constant indep_1 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 77, num_bits );
  constant coef_2 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 97, num_bits );
  constant indep_2 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 467, num_bits );
  constant coef_3 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 286, num_bits );
  constant indep_3 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 1033, num_bits );
  constant coef_4 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 608, num_bits );
  constant indep_4 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 1677, num_bits );
  constant coef_5 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 979, num_bits );
  constant indep_5 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 2048, num_bits );
  constant coef_6 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 608, num_bits );
  constant indep_6 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 2419, num_bits );
  constant coef_7 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 286, num_bits );
  constant indep_7 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 3063, num_bits );
  constant coef_8 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 97, num_bits );
  constant indep_8 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 3629, num_bits );
  constant coef_9 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 10, num_bits );
  constant indep_9 : signed ( ( num_bits - 1 ) downto 0 ) := to_signed( 4019, num_bits );
end package pck_definitions;
